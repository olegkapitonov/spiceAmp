
.subckt 6550_model 1 2 3 4
.param mu=7.9
.param ex=1.35
.param kg1=890
.param kg2=4200
.param kp=60
.param kvb=24
.param  rgi=1000
.param vct=0.0
.param  ccg=14p
.param  cpg1=0.85p
.param  ccp=12p
re1  7 0  1G
e1   7 0  value={v(4,3)/kp*log(1+exp((1/mu+v(2,3)/sqrt(kvb+v(4,3)*v(4,3)))*kp))}
b1   1 3  I='max(pwr(v(7),ex)/kg1*atan(v(1,3)/kvb),0)'
b2   4 3  I='max(pwr(v(4,3)/mu+v(2,3),ex)/kg2,0)'
rcp  1 3  1G
c1   2 3  {ccg}
c2   1 2  {cpg1}
c3   1 3  {ccp}
r1   2 5  {rgi}
d3   5 3  dx
.model dx d(is=1n rs=1 cjo=10pf tt=1n)
.ends
