
.subckt 12AX7_model 1 6 3
.param mu=100
.param ex=1.4
.param kg1=1060
.param kp=600
.param kvb=300
.param  rgi=2000
.param vct=.02
.param  ccg=2.3p
.param  cgp=2.4p
.param  ccp=0.9p
e1 7 0 value='v(1,3)/kp*log(1+exp(kp*(1/mu+v(2,3)/sqrt(kvb+v(1,3)*v(1,3)))))'
re1 7 0 1g
b1 1 3 I = 'max(pwr(v(7),ex)/kg1, 0)'
rcp 1 3 1g
c1 2 3 {ccg}
c2 1 2 {cgp}
c3 1 3 {ccp}
r1 2 5 {rgi}
v1 5 6 {vct}
d3 6 3 dx
.model dx d(is=1n rs=1 cjo=1pf tt=1n)
.ends
